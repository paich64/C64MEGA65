`define BUILD_DATE "2021-07-01"
